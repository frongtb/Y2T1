// Verilog test fixture created from schematic C:\Users\folnw\lab66\lab66.sch - Mon Sep 20 21:44:07 2021

`timescale 1ns / 1ps

module lab66_lab66_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   lab66 UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
